module CSCE611_regfile_testbench;

	logic clk;
	logic rst;
	logic enable;
	logic [15:0] top, next;
	logic [15:0] top_exp, next_exp;
	logic [3:0 ] key;
	logic [1:0 ] mode;
	logic [15:0] val;
	logic [7:0 ] count;

	logic [55:0] vectors [79:0]; 
	logic [55:0] current;
	logic [6:0] i; 

	always begin
		clk = 1'b1; #5;
		clk = 1'b0; #5;
	end
	
	assign rst=({mode,key} == 6'b11_1101) ? 1'b1 : 1'b0;

	rpncalc rpn(.clk(clk),
			.rst(rst),
			.mode(mode),
			.key(key),
			.val(val),
			.top(top),
			.next(next),
			.counter(count));

	initial begin
		// load test vectors from disk
		$readmemh("vectors.dat",vectors);

		for (i = 0; i < 100; i = i + 1) begin

			current = vectors[i];
			
			enable = current[55:55];
			mode = current[53:52];
			key = current[51:48];
			val = current[47:32];
			top_exp = current[31:16];
			next_exp = current[15:0];
			#50;

			if(enable) begin
				$display("current %h",current);
				if (top != top_exp) begin
					$display("Error Top %h", top);
					$display("Top Expected %h",top_exp);
				end
				if (next != next_exp) begin
					$display("Error Next %h", next);
					$display("Next Expected %h",next_exp);
				end
			end

		end 

		// tell the simulator we're done
		$stop();

	end // initial begin

endmodule
