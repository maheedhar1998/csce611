module CSCE611_ri_testbench;
	
endmodule 